��  CCircuit��  CSerializeHack           ��  CPart              ��� 	 CLogicOut�� 	 CTerminal  ����               �            ����           ��    ��  COR
�  `�u�               �          
�  `�u�               �          
�  ����               �            t���           ��    ��  CAND
�  ����                          
�  ����                          
�  ����               �            �|��           ��    �� 	 CInverter
�  � pq                          
�  $p9q              @            d$|           ��    �
�  �  �                           
�   )              @            � �           ��    �
�  � P� Q                          
�  P)Q              @            � D\           ��    ��  CLogicIn�� 	 CLatchKey  X Ah O      !   
�  t H� I                            l Dt L     $    ����     �
�   ��               �          
�   ��     	          �          
�  ,�A�               �            �,�     &      ��    �
�  8�M�               �          
�  8�M�                          
�  d�y�               �            L�d�     *      ��    �
�  8�M�               �          
�  8�M�              @          
�  d�y�     	          �            L�d�     .      ��    �
�  PHeI               �          
�  PXeY              @          
�  |P�Q               �            dD|\     2      ��    �
�  ����              @          
�  ����                          
�  ����               �            ����     6      ��    �
�  �P�Q                          
�  �`�a              @          
�  �X�Y               �            �L�d     :      ��    �
�  � �� �                          
�  �)�              @            � ��     >      ��     �"�  8 yH �      @   
�  T �i �                            L |T �     B    ����      �"�    � 0 �       C   
�  < � Q �                             4 � < �      E    ����                   ���  CWire  ����      G�  x�a�      G�  `�a�       G�  @�a�      G�  x��     	 G�  x�y�      	 G�   x�       G�  �xy      G�  �P�y       G�  �P�Q      G��� 
 CCrossOver  � �         � �      G�S�  � �         � �       G�S�  � D� L        � � �       G�  � ���      G�S�  � D� L        � H� I      G�S�  � �       S�  � l� t        �  � �       G�S�  � L� T        � P� Q      G�  x P� Q      G�  � P�        G�  ���       G�S�  � �         � �� I       G�  �  �       G�  �  �       G�S�  � l� t        � p� q      G�  � ���      G�  � H� I      G�  � H� q       G�  � � q�       G�  P � � �       G�S�  � L� T      S�  � �� �        � � �        G�S�  � �� �        � �� �      G�  � H� �       G�  � �� �       G�  h �y �      G�  x Py �       G�  � �9�      G�  ����       G�  ��	�      G�  �	�       G�  �9�      G�  8pQq      G�  P0Qq       G�  P0!1      G�   �!1       G�   �9�      G�  ���      G�   �9�      G�   ��       G�  P���      G�  P�Q       G�  ( Q      G�   XQY      G�   X!�       G�  (�!�      G�  HQI      G�  H	Y       G�  �X	Y      G�  �`�i       G�  Hh�i      G�  pP�Q      G�  HPIi       G�  (PIQ      G�  p� qQ                     �                             H   K   J    H  j   Y    y  h    }  f    �  _    � $ $ t & N & ' L ' ( ( K * | * + x + , , I . � . / � / 0 0 M 2 � 2 3 � 3 4 4 Q 6 � 6 7 c 7 8 8 � : � : ; � ; < < � > u > ? ? � B B v E E n   , J  I (  M ' L 0 O & P N Q O 4 P R ] U c U e b W W [ R Y W  Z X k l \ T \ i f j _ p a  w b _ U 7 R d V r Z g  o \ h ^ l  \  $ d Z h n � E o o ` o s m g r q d u k x > r B w a v t + z  y { z | { *  ~  } ~ � �  � / 8 � � . � � � 6 � �  � � 3 � � ? � � 2 � � < � ; � � � � : � �  � m �             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 